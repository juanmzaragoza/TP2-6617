----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date: 06/20/2019 12:15:39 PM
-- Design Name: 
-- Module Name: font_ROM - Behavioral
-- Project Name: 
-- Target Devices: 
-- Tool Versions: 
-- Description: 
-- 
-- Dependencies: 
-- 
-- Revision:
-- Revision 0.01 - File Created
-- Additional Comments:
-- 
----------------------------------------------------------------------------------


library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx leaf cells in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

-- TODO: la idea es que los caracteres sean de 8x8 (2^3x8)
-- en este caso, tenemos caracters de 16x8 (2^4x8) => REDUCIR!
--
-- Los primeros 7 bits de addrA nos van a devolver el caracter
-- mientras que los ultimos AW-7 bits nos van a devolver los
-- 8 bits correspondientes a la fila del caracter
entity font_ROM is
    generic(
		AW: integer := 11; -- usar 2^10
		DW: integer := 8
	);
	port(
		--clkA: in std_logic;
		--writeEnableA: in std_logic := '0'; -- NO USAR
		addrIn: in std_logic_vector(AW-1 downto 0);
		--dataInA: in std_logic_vector(DW-1 downto 0) := (others => '0'); -- NO USAR
		dataOut: out std_logic_vector(DW-1 downto 0)
	);
end font_ROM;

architecture Behavioral of font_ROM is



	type rom_type is array (0 to 2**AW-1) of std_logic_vector(DW-1 downto 0);

	-- ROM definition
	signal ROM: rom_type := (   -- 2^11-by-8
		-- NUL: code x00
		"00000000", -- 0
		"00000000", -- 1
		"00000000", -- 2
		"00000000", -- 3
		"00000000", -- 4
		"00000000", -- 5
		"00000000", -- 6
		"00000000", -- 7
		-- SOH: code x01
		"01111110", -- 0  ******
		"10000001", -- 1 *      *
		"10100101", -- 2 * *  * *
		"10000001", -- 3 *      *
		"10111101", -- 4 * **** *
		"10011001", -- 5 *  **  *
		"10000001", -- 6 *      *
		"01111110", -- 7  ******
		-- STX: code x02
		"01111110", -- 0  ******
		"11111111", -- 1 ********
		"11011011", -- 2 ** ** **
		"11111111", -- 3 ********
		"11000011", -- 4 **    **
		"11100111", -- 5 ***  ***
		"11111111", -- 6 ********
		"01111110", -- 7  ******
		-- ETX: code x03
		"01101100", -- 4  ** **
		"11111110", -- 5 *******
		"11111110", -- 6 *******
		"11111110", -- 7 *******
		"11111110", -- 8 *******
		"01111100", -- 9  *****
		"00111000", -- a   ***
		"00010000", -- b    *
		-- EOT: code x04
		"00000000", -- 0
		"00010000", -- 1    *
		"00111000", -- 2   ***
		"01111100", -- 3  *****
		"11111110", -- 4 *******
		"01111100", -- 5  *****
		"00111000", -- 6   ***
		"00010000", -- 7    *
		-- ENQ: code x05
		"00011000", -- 3    **
		"00111100", -- 5   ****
		"11100111", -- 6 ***  ***
		"11100111", -- 7 ***  ***
		"11100111", -- 8 ***  ***
		"00011000", -- 9    **
		"00011000", -- a    **
		"00111100", -- b   ****
		-- ACK: code x06
		"00011000", -- 3    **
		"00111100", -- 4   ****
		"01111110", -- 5  ******
		"11111111", -- 6 ********
		"01111110", -- 8  ******
		"00011000", -- 9    **
		"00011000", -- a    **
		"00111100", -- b   ****
		-- BEL: code x07
		"00000000", -- 0
		"00000000", -- 1
		"00000000", -- 2
		"00000000", -- 3
		"00011000", -- 4    **
		"00111100", -- 5   ****
		"00111100", -- 6   ****
		"00011000", -- 7    **
		-- BS: code x08
		"11111111", -- 0 ********
		"11111111", -- 1 ********
		"11100111", -- 2 ***  ***
		"11000011", -- 3 **    **
		"11000011", -- 4 **    **
		"11100111", -- 5 ***  ***
		"11111111", -- 6 ********
		"11111111", -- 7 ********
		-- HT: code x09
		"00000000", -- 0
		"00000000", -- 1
		"00111100", -- 2   ****
		"01100110", -- 3  **  **
		"01000010", -- 4  *    *
		"01000010", -- 5  *    *
		"01100110", -- 6  **  **
		"00111100", -- 7   ****
		-- LF: code x0a
		"11111111", -- 0 ********
		"11000011", -- 1 **    **
		"10011001", -- 2 *  **  *
		"10111101", -- 3 * **** *
		"10111101", -- 4 * **** *
		"10011001", -- 5 *  **  *
		"11000011", -- 6 **    **
		"11111111", -- 7 ********
		-- code x0b
		"00011110", -- 0    ****
		"00001110", -- 1     ***
		"00011010", -- 2    ** *
		"00110010", -- 3   **  *
		"01111000", -- 4  ****
		"11001100", -- 5 **  **
		"11001100", -- 6 **  **
		"01111000", -- 7  ****
		-- code x0c
		"00111100", -- 0   ****
		"01100110", -- 1  **  **
		"01100110", -- 2  **  **
		"00111100", -- 3   ****
		"00011000", -- 4    **
		"01111110", -- 5  ******
		"00011000", -- 6    **
		"00011000", -- 7    **
		-- code x0d
		"00111111", -- 0   ******
		"00110011", -- 1   **  **
		"00111111", -- 2   ******
		"00110000", -- 3   **
		"00110000", -- 4   **
		"01110000", -- 5  ***
		"11110000", -- 6 ****
		"11100000", -- 7 ***
		-- code x0e
		"01111111", -- 0  *******
		"01100011", -- 1  **   **
		"01111111", -- 2  *******
		"01100011", -- 3  **   **
		"01100111", -- 4  **  ***
		"11100111", -- 5 ***  ***
		"11100110", -- 6 ***  **
		"11000000", -- 7 **
		-- code x0f
		"00011000", -- 0    **
		"11011011", -- 1 ** ** **
		"00111100", -- 2   ****
		"11100111", -- 3 ***  ***
		"00111100", -- 4   ****
		"11011011", -- 5 ** ** **
		"00011000", -- 6    **
		"00011000", -- 7    **
		-- code x10
		"10000000", -- 0 *
		"11000000", -- 1 **
		"11100000", -- 2 ***
		"11110000", -- 3 ****
		"11111000", -- 4 *****
		"11110000", -- 5 ****
		"11100000", -- 6 ***
		"11000000", -- 7 **
		-- code x11
		"00000010", -- 0       *
		"00000110", -- 1      **
		"00001110", -- 2     ***
		"00011110", -- 3    ****
		"00111110", -- 4   *****
		"00011110", -- 5    ****
		"00001110", -- 6     ***
		"00000110", -- 7      **
		-- code x12
		"00011000", -- 0    **
		"00111100", -- 1   ****
		"01111110", -- 2  ******
		"00011000", -- 3    **
		"00011000", -- 4    **
		"01111110", -- 5  ******
		"00111100", -- 6   ****
		"00011000", -- 7    **
		-- code x13
		"01100110", -- 0  **  **
		"01100110", -- 1  **  **
		"01100110", -- 2  **  **
		"01100110", -- 3  **  **
		"01100110", -- 4  **  **
		"00000000", -- 5
		"01100110", -- 6  **  **
		"01100110", -- 7  **  **
		-- code x14
		"01111111", -- 0  *******
		"11011011", -- 1 ** ** **
		"11011011", -- 2 ** ** **
		"11011011", -- 3 ** ** **
		"01111011", -- 4  **** **
		"00011011", -- 5    ** **
		"00011011", -- 6    ** **
		"00011011", -- 7    ** **
		-- code x15
		"01111100", -- 0  *****
		"11000110", -- 1 **   **
		"01100000", -- 2  **
		"01101100", -- 3  ** **
		"01101100", -- 4  ** **
		"00001100", -- 5     **
		"11000110", -- 6 **   **
		"01111100", -- 7  *****
		-- code x16
		"00000000", -- 0
		"00000000", -- 1
		"00000000", -- 2
		"00000000", -- 3
		"11111110", -- 4 *******
		"11111110", -- 5 *******
		"11111110", -- 6 *******
		"11111110", -- 7 *******
		-- code x17
		"00011000", -- 0    **
		"00111100", -- 1   ****
		"01111110", -- 2  ******
		"00011000", -- 3    **
		"01111110", -- 4  ******
		"00111100", -- 5   ****
		"00011000", -- 6    **
		"01111110", -- 7  ******
		-- code x18
		"00011000", -- 0    **
		"00111100", -- 1   ****
		"01111110", -- 2  ******
		"00011000", -- 3    **
		"00011000", -- 4    **
		"00011000", -- 5    **
		"00011000", -- 6    **
		"00011000", -- 7    **
		-- code x19
		"00011000", -- 0    **
		"00011000", -- 1    **
		"00011000", -- 2    **
		"00011000", -- 3    **
		"00011000", -- 4    **
		"01111110", -- 5  ******
		"00111100", -- 6   ****
		"00011000", -- 7    **
		-- code x1a
		"00000000", -- 0
		"00000000", -- 1
		"00000000", -- 2
		"00011000", -- 3    **
		"00001100", -- 4     **
		"11111110", -- 5 *******
		"00001100", -- 6     **
		"00011000", -- 7    **
		-- code x1b
		"00000000", -- 0
		"00000000", -- 1
		"00000000", -- 2
		"00110000", -- 3   **
		"01100000", -- 4  **
		"11111110", -- 5 *******
		"01100000", -- 6  **
		"00110000", -- 7   **
		-- code x1c
		"00000000", -- 0
		"00000000", -- 1
		"00000000", -- 2
		"00000000", -- 3
		"11000000", -- 4 **
		"11000000", -- 5 **
		"11000000", -- 6 **
		"11111110", -- 7 *******
		-- code x1d
		"00000000", -- 0
		"00000000", -- 1
		"00000000", -- 2
		"00100100", -- 3   *  *
		"01100110", -- 4  **  **
		"11111111", -- 5 ********
		"01100110", -- 6  **  **
		"00100100", -- 7   *  *
		-- code x1e
		"00000000", -- 0
		"00010000", -- 1    *
		"00111000", -- 2   ***
		"00111000", -- 3   ***
		"01111100", -- 4  *****
		"01111100", -- 5  *****
		"11111110", -- 6 *******
		"11111110", -- 7 *******
		-- code x1f
		"00000000", -- 0
		"11111110", -- 1 *******
		"11111110", -- 2 *******
		"01111100", -- 3  *****
		"01111100", -- 4  *****
		"00111000", -- 5   ***
		"00111000", -- 6   ***
		"00010000", -- 7    *
		-- code x20
		"00000000", -- 0
		"00000000", -- 1
		"00000000", -- 2
		"00000000", -- 3
		"00000000", -- 4
		"00000000", -- 5
		"00000000", -- 6
		"00000000", -- 7
		-- code x21
		"00011000", -- 0    **
		"00111100", -- 1   ****
		"00111100", -- 2   ****
		"00011000", -- 3    **
		"00011000", -- 4    **
		"00000000", -- 5
		"00011000", -- 6    **
		"00011000", -- 7    **
		-- code x22
		"00000000", -- 0
		"01100110", -- 1  **  **
		"01100110", -- 2  **  **
		"01100110", -- 3  **  **
		"00100100", -- 4   *  *
		"00000000", -- 5
		"00000000", -- 6
		"00000000", -- 7
		-- code x23
		"01101100", -- 0  ** **
		"01101100", -- 1  ** **
		"11111110", -- 2 *******
		"01101100", -- 3  ** **
		"01101100", -- 4  ** **
		"11111110", -- 5 *******
		"01101100", -- 6  ** **
		"01101100", -- 7  ** **
		-- code x24
		"00111000", -- 0    ***
		"11000010", -- 1  **    *
		"11000000", -- 2  **
		"01111100", -- 3   *****
		"00000110", -- 4       **
		"10000110", -- 5  *    **
		"01111100", -- 6   *****
		"00011000", -- 7     **
		-- code x25
		"11000010", -- 0 **    *
		"11000110", -- 1 **   **
		"00001100", -- 2     **
		"00011000", -- 3    **
		"00110000", -- 4   **
		"01100000", -- 5  **
		"11000110", -- 6 **   **
		"10000110", -- 7 *    **
		-- code x26
		"00111000", -- 0   ***
		"01101100", -- 1  ** **
		"01101100", -- 2  ** **
		"00111000", -- 3   ***
		"01110110", -- 4  *** **
		"11011100", -- 5 ** ***
		"11001100", -- 6 **  **
		"01110110", -- 7  *** **
		-- code x27
		"00000000", -- 0
		"00110000", -- 1   **
		"00110000", -- 2   **
		"00110000", -- 3   **
		"01100000", -- 4  **
		"00000000", -- 5
		"00000000", -- 6
		"00000000", -- 7
		-- code x28
		"00001100", -- 0     **
		"00011000", -- 1    **
		"00110000", -- 2   **
		"00110000", -- 3   **
		"00110000", -- 4   **
		"00110000", -- 5   **
		"00011000", -- 6    **
		"00001100", -- 7     **
		-- code x29
		"00110000", -- 0   **
		"00011000", -- 1    **
		"00001100", -- 2     **
		"00001100", -- 3     **
		"00001100", -- 4     **
		"00001100", -- 5     **
		"00011000", -- 6    **
		"00110000", -- 7   **
		-- code x2a
		"00000000", -- 0
		"00000000", -- 1
		"00000000", -- 2
		"01100110", -- 3  **  **
		"00111100", -- 4   ****
		"11111111", -- 5 ********
		"00111100", -- 6   ****
		"01100110", -- 7  **  **
		-- code x2b
		"00000000", -- 0
		"00000000", -- 1
		"00000000", -- 2
		"00011000", -- 3    **
		"00011000", -- 4    **
		"01111110", -- 5  ******
		"00011000", -- 6    **
		"00011000", -- 7    **
		-- code x2c
		"00000000", -- 0
		"00000000", -- 1
		"00000000", -- 2
		"00000000", -- 3
		"00011000", -- 4    **
		"00011000", -- 5    **
		"00011000", -- 6    **
		"00110000", -- 7   **
		-- code x2d
		"00000000", -- 0
		"00000000", -- 1
		"00000000", -- 2
		"00000000", -- 3
		"01111110", -- 4  ******
		"00000000", -- 5
		"00000000", -- 6
		"00000000", -- 7
		-- code x2e
		"00000000", -- 0
		"00000000", -- 1
		"00000000", -- 2
		"00011000", -- 3    **
		"00011000", -- 4    **
		"00000000", -- 5
		"00000000", -- 6
		"00000000", -- 7
		-- code x2f
		"00000010", -- 0       *
		"00000110", -- 1      **
		"00001100", -- 2     **
		"00011000", -- 3    **
		"00110000", -- 4   **
		"01100000", -- 5  **
		"11000000", -- 6 **
		"10000000", -- 7 *
		-- 0: code x30
		"01111100", -- 0  *****
		"11000110", -- 1 **   **
		"11001110", -- 2 **  ***
		"11011110", -- 3 ** ****
		"11110110", -- 4 **** **
		"11100110", -- 5 ***  **
		"11000110", -- 6 **   **
		"01111100", -- 7  *****
		-- 1: code x31
		"01111000", -- 0    **
		"00011000", -- 1   ***
		"00011000", -- 2  ****
		"00011000", -- 3    **
		"00011000", -- 4    **
		"00011000", -- 5    **
		"00011000", -- 6    **
		"01111110", -- 7  ******
		-- 2: code x32
		"01111100", -- 0  *****
		"11000110", -- 1 **   **
		"00001100", -- 2     **
		"00011000", -- 3    **
		"00110000", -- 4   **
		"01100000", -- 5  **
		"11000110", -- 6 **   **
		"11111110", -- 7 *******
		-- 3: code x33
		"01111100", -- 0  *****
		"11000110", -- 1 **   **
		"00000110", -- 2      **
		"00111100", -- 3   ****
		"00000110", -- 4      **
		"00000110", -- 5      **
		"11000110", -- 6 **   **
		"01111100", -- 7  *****
		-- 4: code x34
		"00001100", -- 0     **
		"00011100", -- 1    ***
		"01101100", -- 2  ** **
		"11001100", -- 3 **  **
		"11111110", -- 4 *******
		"00001100", -- 5     **
		"00001100", -- 6     **
		"00011110", -- 7    ****
		-- code x35
		"11111110", -- 0 *******
		"11000000", -- 1 **
		"11000000", -- 2 **
		"11111100", -- 3 ******
		"00000110", -- 4      **
		"00000110", -- 5      **
		"11000110", -- 6 **   **
		"01111100", -- 7  *****
		-- code x36
		"00111000", -- 0   ***
		"01100000", -- 1  **
		"11000000", -- 2 **
		"11000000", -- 3 **
		"11111100", -- 4 ******
		"11000110", -- 5 **   **
		"11000110", -- 6 **   **
		"01111100", -- 7  *****
		-- code x37
		"11111110", -- 0 *******
		"11000110", -- 1 **   **
		"00000110", -- 2      **
		"00001100", -- 3     **
		"00011000", -- 4    **
		"00110000", -- 5   **
		"00110000", -- 6   **
		"00110000", -- 7   **
		-- code x38
		"01111100", -- 0  *****
		"11000110", -- 1 **   **
		"11000110", -- 2 **   **
		"01111100", -- 3  *****
		"11000110", -- 4 **   **
		"11000110", -- 5 **   **
		"11000110", -- 6 **   **
		"01111100", -- 7  *****
		-- code x39
		"01111100", -- 0  *****
		"11000110", -- 1 **   **
		"11000110", -- 2 **   **
		"11000110", -- 3 **   **
		"01111110", -- 4  ******
		"00000110", -- 5      **
		"00001100", -- 6     **
		"01111000", -- 7  ****
		-- code x3a
		"00000000", -- 0
		"00011000", -- 1    **
		"00011000", -- 2    **
		"00000000", -- 3
		"00000000", -- 4
		"00011000", -- 5    **
		"00011000", -- 6    **
		"00000000", -- 7
		-- code x3b=
		"00000000", -- 0
		"00011000", -- 1    **
		"00011000", -- 2    **
		"00000000", -- 3
		"00000000", -- 4
		"00011000", -- 5    **
		"00110000", -- 6   **
		"00000000", -- 7
		-- code x3c
		"00000110", -- 0      **
		"00001100", -- 1     **
		"00011000", -- 2    **
		"00110000", -- 3   **
		"01100000", -- 4  **
		"00110000", -- 5   **
		"00011000", -- 6    **
		"00001100", -- 7     **
		-- code x3d
		"00000000", -- 0
		"00000000", -- 1
		"01111110", -- 2  ******
		"00000000", -- 3
		"00000000", -- 4
		"01111110", -- 5  ******
		"00000000", -- 6
		"00000000", -- 7
		-- code x3e
		"01100000", -- 0  **
		"00110000", -- 1   **
		"00011000", -- 2    **
		"00001100", -- 3     **
		"00000110", -- 4      **
		"00001100", -- 5     **
		"00011000", -- 6    **
		"00110000", -- 7   **
		-- code x3f
		"01111100", -- 0  *****
		"11000110", -- 1 **   **
		"00001100", -- 2     **
		"00011000", -- 3    **
		"00011000", -- 4    **
		"00000000", -- 5
		"00011000", -- 6    **
		"00011000", -- 7    **
		-- code x40
		"01111100", -- 0  *****
		"11000110", -- 1 **   **
		"11000110", -- 2 **   **
		"11011110", -- 3 ** ****
		"11011110", -- 4 ** ****
		"11011100", -- 5 ** ***
		"11000000", -- 6 **
		"01111100", -- 7  *****
-- Tabla de mayusculas ASCII 8x8
	
		-- A: code x41
		
	"01110000", 
	"10001000",
	"10001000",
	"10001000",
	"11111000",
	"10001000",
	"10001000",
	"00000000",
		
		-- B: code x42
	
	"11110000", 
	"10001000",
	"10001000",
	"11110000",
	"10001000",	
	"10001000",
	"11110000",
	"00000000",
		
		-- C: code x43
	
	"01110000", 
	"10001000",
	"10000000",
	"10000000",
	"10000000",	
	"10001000",
	"01110000",
	"00000000",
		
		-- D: code x44
	
	"11110000", 
	"10001000",
	"10001000",
	"10001000",
	"10001000",	
	"10001000",
	"11110000",
	"00000000",
		
		-- E :code x45
	
	"11111000", 
	"10000000",
	"10000000",
	"11100000",
	"10000000",	
	"10000000",
	"11111000",
	"00000000",
		
		-- F: code x46
	
	"11111000", 
	"10000000",
	"10000000",
	"11100000",
	"10000000",	
	"10000000",
	"10000000",
	"00000000",
		
		-- G: code x47
		
	"01110000", 
	"10001000",
	"10000000",
	"10111000",
	"10001000",	
	"10001000",
	"01110000",
	"00000000",
		
		-- H: code x48
	
	"10001000", 
	"10001000",
	"10001000",
	"11111000",
	"10001000",	
	"10001000",
	"10001000",
	"00000000",
		
		-- I: code x49
	
	"01110000", 
	"00100000",
	"00100000",
	"00100000",
	"00100000",	
	"00100000",
	"01110000",
	"00000000",
		
		-- J: code x4a
	
	"00111000", 
	"00010000",
	"00010000",
	"00010000",
	"00010000",	
	"10010000",
	"01100000",
	"00000000",
		
		-- K: code x4b
	
	"10001000", 
	"10010000",
	"10100000",
	"11000000",
	"10100000",	
	"10010000",
	"10001000",
	"00000000",
		
		-- L: code x4c
	
	"10000000", 
	"10000000",
	"10000000",
	"10000000",
	"10000000",	
	"10000000",
	"11111000",
	"00000000",
		
		-- M: code x4d
	
	"10001000", 
	"11011000",
	"10101000",
	"10001000",
	"10001000",	
	"10001000",
	"10001000",
	"00000000",
		
		-- N: code x4e
	
	"10001000", 
	"10001000",
	"11001000",
	"10101000",
	"10011000",	
	"10001000",
	"10001000",
	"00000000",
		
		-- O: code x4f
	
	"01110000", 
	"10001000",
	"10001000",
	"10001000",
	"10001000",	
	"10001000",
	"01110000",
	"00000000",
		
		-- P: code x50
	
	"11110000", 
	"10001000",
	"10001000",
	"11110000",
	"10000000",	
	"10000000",
	"10000000",
	"00000000",
		
		-- Q: code x510
	
	"01110000", 
	"10001000",
	"10001000",
	"10001000",
	"10101000",	
	"10010000",
	"01101000",
	"00000000",
	
		-- R: code x52
	
	"11110000", 
	"10001000",
	"10001000",
	"11110000",
	"10100000",	
	"10010000",
	"10001000",
	"00000000",
		
		-- S: code x53
	
	"01111000", 
	"10000000",
	"10000000",
	"01110000",
	"00001000",	
	"00001000",
	"11110000",
	"00000000",
		
		-- T: code x54
	
	"11111000", 
	"00100000",
	"00100000",
	"00100000",
	"00100000",	
	"00100000",
	"00100000",
	"00000000",
		
		-- U: code x55
	
	"10001000", 
	"10001000",
	"10001000",
	"10001000",
	"10001000",	
	"10001000",
	"01110000",
	"00000000",
		
		-- V: code x56
	
	"10001000", 
	"10001000",
	"10001000",
	"10001000",
	"10001000",	
	"01010000",
	"00100000",
	"00000000",		
		-- W: code x57
	
	"10001000", 
	"10001000",
	"10001000",
	"10001000",
	"10101000",	
	"10101000",
	"01010000",
	"00000000",
		

		-- X: code x58
	
	"10001000", 
	"10001000",
	"01010000",
	"00100000",
	"01010000",	
	"10001000",
	"10001000",
	"00000000",
		
		-- Y: code x59
	
	"10001000", 
	"10001000",
	"10001000",
	"01010000",
	"00100000",	
	"00100000",
	"00100000",
	"00000000",
	

		
		-- Z: code x5a
	
	"11111000", 
	"00001000",
	"00010000",
	"00100000",
	"01000000",	
	"10000000",
	"11111000",
	"00000000",
		
		
		-- code x5b
		"00111100", -- 0   ****
		"00110000", -- 1   **
		"00110000", -- 2   **
		"00110000", -- 3   **
		"00110000", -- 4   **
		"00110000", -- 5   **
		"00110000", -- 6   **
		"00111100", -- 7   ****
		-- code x5c
		"10000000", -- 0 *
		"11000000", -- 1 **
		"11100000", -- 2 ***
		"01110000", -- 3  ***
		"00111000", -- 4   ***
		"00001110", -- 5     ***
		"00000110", -- 6      **
		"00000010", -- 7       *
		-- code x5d
		"00111100", -- 0   ****
		"00001100", -- 1     **
		"00001100", -- 2     **
		"00001100", -- 3     **
		"00001100", -- 4     **
		"00001100", -- 5     **
		"00001100", -- 6     **
		"00111100", -- 7   ****
		-- code x5e
		"00010000", -- 0    *
		"00111000", -- 1   ***
		"01101100", -- 2  ** **
		"11000110", -- 3 **   **
		"00000000", -- 4
		"00000000", -- 5
		"00000000", -- 6
		"00000000", -- 7
		-- code x5f
		"00000000", -- 0
		"00000000", -- 1
		"00000000", -- 2
		"00000000", -- 3
		"00000000", -- 4
		"11111111", -- 5 ********
		"00000000", -- 6
		"00000000", -- 7
		-- code x60
		"00110000", -- 0   **
		"00110000", -- 1   **
		"00011000", -- 2    **
		"00000000", -- 3
		"00000000", -- 4
		"00000000", -- 5
		"00000000", -- 6
		"00000000", -- 7
		-- a: code x61
		"00000000", -- 0
		"01111000", -- 1  ****
		"00001100", -- 2     **
		"01111100", -- 3  *****
		"11001100", -- 4 **  **
		"11001100", -- 5 **  **
		"11001100", -- 6 **  **
		"01110110", -- 7  *** **
		-- b: code x62
		"00000000", -- 0
		"11100000", -- 1  ***
		"01100000", -- 2   **
		"01100000", -- 3   **
		"01111000", -- 4   ****
		"01101100", -- 5   ** **
		"01100110", -- 6   **  **
		"01111100", -- 7   *****
		-- c: code x63
		"00000000", -- 0
		"00000000", -- 1
		"01111100", -- 2  *****
		"11000110", -- 3 **   **
		"11000000", -- 4 **
		"11000000", -- 5 **
		"11000110", -- 6 **   **
		"01111100", -- 7  *****
		-- d: code x64
		"00000000", -- 0
		"00000000", -- 1
		"00011100", -- 2    ***
		"00001100", -- 3     **
		"00111100", -- 4   ****
		"01101100", -- 5  ** **
		"11001100", -- 6 **  **
		"01110110", -- 7  *** **
		-- e: code x65
		"00000000", -- 0
		"01111100", -- 1  *****
		"11000110", -- 2 **   **
		"11111110", -- 3 *******
		"11000000", -- 4 **
		"11000000", -- 5 **
		"11000110", -- 6 **   **
		"01111100", -- 7  *****
		-- f: code x66
		"00000000", -- 0
		"00111000", -- 1   ***
		"01100100", -- 2  **  *
		"01100000", -- 3  **
		"11110000", -- 4 ****
		"01100000", -- 5  **
		"01100000", -- 6  **
		"11110000", -- 7 ****
		-- g: code x67
		"00000000", -- 0
		"01110110", -- 1  *** **
		"11001100", -- 2 **  **
		"11001100", -- 3 **  **
		"01111100", -- 4  *****
		"00001100", -- 5     **
		"11001100", -- 6 **  **
		"01111000", -- 7  ****
		-- h: code x68
		"00000000", -- 0
		"11100000", -- 1 ***
		"01100000", -- 2  **
		"01100000", -- 3  **
		"01101100", -- 4  ** **
		"01110110", -- 5  *** **
		"01100110", -- 6  **  **
		"11100110", -- 7 ***  **
		-- i: code x69
		"00000000", -- 0
		"00011000", -- 1    **
		"00011000", -- 2    **
		"00000000", -- 3
		"00111000", -- 4   ***
		"00011000", -- 5    **
		"00011000", -- 6    **
		"00111100", -- 7   ****
		-- j: code x6a
		"00000000", -- 0
		"00000110", -- 1      **
		"00000110", -- 2      **
		"00000000", -- 3
		"00001110", -- 4     ***
		"00000110", -- 5      **
		"01100110", -- 6  **  **
		"00111100", -- 7   ****
		-- k: code x6b
		"11100000", -- 0 ***
		"01100000", -- 1  **
		"01100110", -- 2  **  **
		"01101100", -- 3  ** **
		"01111000", -- 4  ****
		"01101100", -- 5  ** **
		"01100110", -- 6  **  **
		"11100110", -- 7 ***  **
		-- l: code x6c
		"00000000", -- 0
		"00111000", -- 1   ***
		"00011000", -- 2    **
		"00011000", -- 3    **
		"00011000", -- 4    **
		"00011000", -- 5    **
		"00011000", -- 6    **
		"00111100", -- 7   ****
		-- m: code x6d
		"00000000", -- 0
		"11100110", -- 1 ***  **
		"11111111", -- 2 ********
		"11011011", -- 3 ** ** **
		"11011011", -- 4 ** ** **
		"11011011", -- 5 ** ** **
		"11011011", -- 6 ** ** **
		"11011011", -- 7 ** ** **
		-- n: code x6e
		"00000000", -- 0
		"11011100", -- 1 ** ***
		"01100110", -- 2  **  **
		"01100110", -- 3  **  **
		"01100110", -- 4  **  **
		"01100110", -- 5  **  **
		"01100110", -- 6  **  **
		"01100110", -- 7  **  **
		-- o: code x6f
		"00000000", -- 0
		"01111100", -- 1  *****
		"11000110", -- 2 **   **
		"11000110", -- 3 **   **
		"11000110", -- 4 **   **
		"11000110", -- 5 **   **
		"11000110", -- 6 **   **
		"01111100", -- 7  *****
		-- code x70
		"00000000", -- 0
		"11011100", -- 1 ** ***
		"01100110", -- 2  **  **
		"01100110", -- 3  **  **
		"01111100", -- 4  *****
		"01100000", -- 5  **
		"01100000", -- 6  **
		"11110000", -- 7 ****
		-- code x71
		"00000000", -- 0
		"01110110", -- 1  *** **
		"11001100", -- 2 **  **
		"11001100", -- 3 **  **
		"11001100", -- 4 **  **
		"01111100", -- 5  *****
		"00001100", -- 6     **
		"00011110", -- 7    ****
		-- code x72
		"00000000", -- 0
		"11011100", -- 1 ** ***
		"01110110", -- 2  *** **
		"01100110", -- 3  **  **
		"01100000", -- 4  **
		"01100000", -- 5  **
		"01100000", -- 6  **
		"11110000", -- 7 ****
		-- code x73
		"00000000", -- 0
		"01111100", -- 1  *****
		"11000110", -- 2 **   **
		"01100000", -- 3  **
		"00111000", -- 4   ***
		"00001100", -- 5     **
		"11000110", -- 6 **   **
		"01111100", -- 7  *****
		-- code x74
		"00000000", -- 0
		"00010000", -- 1    *
		"00110000", -- 2   **
		"11111100", -- 3 ******
		"00110000", -- 4   **
		"00110000", -- 5   **
		"00110110", -- 6   ** **
		"00011100", -- 7    ***
		-- code x75
		"00000000", -- 0
		"11001100", -- 1 **  **
		"11001100", -- 2 **  **
		"11001100", -- 3 **  **
		"11001100", -- 4 **  **
		"11001100", -- 5 **  **
		"11001100", -- 6 **  **
		"01110110", -- 7  *** **
		-- code x76
		"00000000", -- 0
		"11000011", -- 1 **    **
		"11000011", -- 2 **    **
		"11000011", -- 3 **    **
		"11000011", -- 4 **    **
		"01100110", -- 5  **  **
		"00111100", -- 6   ****
		"00011000", -- 7    **
		-- code x77
		"00000000", -- 0
		"11000011", -- 1 **    **
		"11000011", -- 2 **    **
		"11000011", -- 3 **    **
		"11011011", -- 4 ** ** **
		"11011011", -- 5 ** ** **
		"11111111", -- 6 ********
		"01100110", -- 7  **  **
		-- code x78
		"00000000", -- 0
		"11000011", -- 1 **    **
		"01100110", -- 2  **  **
		"00111100", -- 3   ****
		"00011000", -- 4    **
		"00111100", -- 5   ****
		"01100110", -- 6  **  **
		"11000011", -- 7 **    **
		-- code x79
		"00000000", -- 0
		"11000110", -- 1 **   **
		"11000110", -- 2 **   **
		"11000110", -- 3 **   **
		"01111110", -- 4  ******
		"00000110", -- 5      **
		"00001100", -- 6     **
		"11111000", -- 7 *****
		-- code x7a
		"00000000", -- 0
		"11111110", -- 1 *******
		"11001100", -- 2 **  **
		"00011000", -- 3    **
		"00110000", -- 4   **
		"01100000", -- 5  **
		"11000110", -- 6 **   **
		"11111110", -- 7 *******
		-- code x7b
		"00001110", -- 0     ***
		"00011000", -- 1    **
		"00011000", -- 2    **
		"01110000", -- 3  ***
		"00011000", -- 4    **
		"00011000", -- 5    **
		"00011000", -- 6    **
		"00001110", -- 7     ***
		-- code x7c
		"00011000", -- 0    **
		"00011000", -- 1    **
		"00011000", -- 2    **
		"00000000", -- 3
		"00011000", -- 4    **
		"00011000", -- 5    **
		"00011000", -- 6    **
		"00011000", -- 7    **
		-- code x7d
		"01110000", -- 0  ***
		"00011000", -- 1    **
		"00011000", -- 2    **
		"00001110", -- 3     ***
		"00011000", -- 4    **
		"00011000", -- 5    **
		"00011000", -- 6    **
		"01110000", -- 7  ***
		-- code x7e
		"01110110", -- 0  *** **
		"11011100", -- 1 ** ***
		"00000000", -- 2
		"00000000", -- 3
		"00000000", -- 4
		"00000000", -- 5
		"00000000", -- 6
		"00000000", -- 7
		-- code x7f
		"00010000", -- 0    *
		"00111000", -- 1   ***
		"01101100", -- 2  ** **
		"11000110", -- 3 **   **
		"11000110", -- 4 **   **
		"11000110", -- 5 **   **
		"11111110", -- 6 *******
		"00000000"  -- 7
	);
	
begin

	-- addr register to infer block RAM
--	setRegA: process (clkA)
--	begin
--		if rising_edge(clkA) then
		
--			-- Write to rom
--			if(writeEnableA = '1') then
--				ROM(to_integer(unsigned(addrA))) <= dataInA;
--			end if;

--		end if;
--	end process;
    
    -- Read from it
    dataOut <= ROM(to_integer(unsigned(addrIn)));

end Behavioral;
